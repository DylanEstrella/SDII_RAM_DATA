--32-word 8-bit synchronous RAM with enable
--https://github.com/VHDL-Digital-Systems
--http://blog.espol.edu.ec/sistemasdigitalesfiec

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ram_type_pck is
	type ram_type is array (0 to (2**8)-1) of std_logic_vector(8-1 downto 0);
end package;



--Library
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.ram_type_pck.all;

--Entity
entity SRAM is 
	generic(n: integer:=8;-- n-bits per data
	m: integer:=8); -- m-bits of addresses
	port(
		clk,en,wr: in std_logic;
		info: in ram_type;
		addr : in std_logic_vector(m-1 downto 0); 
		Din : in std_logic_vector(n-1 downto 0);
		Dout : out std_logic_vector(n-1 downto 0)); 
end SRAM;

--Architecture
architecture solve of SRAM is
	-- Signals,Constants,Variables,Components	
	--type ram_type is array (0 to (2**m)-1) of std_logic_vector(n-1 downto 0); 
	signal tmp_ram: ram_type:=(
		b"00000011",
		b"00000100",
		b"00000101",
		b"00000110",
		b"00000111",
		b"00001000",
		b"00001001",
		b"00001010",
		b"00001011",
		b"00001100",
		b"00001101",
		b"00001110",
		b"00001111",
		b"00010000",
		b"00010001",
		b"00010010",
		b"00010011",
		b"00010100",
		b"00010101",
		b"00010110",
		b"00010111",
		b"00011000",
		b"00011001",
		b"00011010",
		b"00011011",
		b"00011100",
		b"00011101",
		b"00011110",
		b"00011111",
		b"00100000",
		b"00100001",
		b"00100010",
		b"00100011",
		b"00100100",
		b"00100101",
		b"00100110",
		b"00100111",
		b"00101000",
		b"00101001",
		b"00101010",
		b"00101011",
		b"00101100",
		b"00101101",
		b"00101110",
		b"00101111",
		b"00110000",
		b"00110001",
		b"00110010",
		b"00110011",
		b"00110100",
		b"00110101",
		b"00110110",
		b"00110111",
		b"00111000",
		b"00111001",
		b"00111010",
		b"00111011",
		b"00111100",
		b"00111101",
		b"00111110",
		b"00111111",
		b"01000000",
		b"01000001",
		b"01000010",
		b"01000011",
		b"01000100",
		b"01000101",
		b"01000110",
		b"01000111",
		b"01001000",
		b"01001001",
		b"01001010",
		b"01001011",
		b"01001100",
		b"01001101",
		b"01001110",
		b"01001111",
		b"01010000",
		b"01010001",
		b"01010010",
		b"01010011",
		b"01010100",
		b"01010101",
		b"01010110",
		b"01010111",
		b"01011000",
		b"01011001",
		b"01011010",
		b"01011011",
		b"01011100",
		b"01011101",
		b"01011110",
		b"01011111",
		b"01100000",
		b"01100001",
		b"01100010",
		b"01100011",
		b"01100100",
		b"01100101",
		b"01100110",
		b"01100111",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000",
		b"00000000",b"00000000",b"00000000",b"00000000",b"00000000"
	 ); 
	begin
	--Process #1:
	process(clk,wr)
	--Sequential programming
		begin
			if (clk'event and clk='1') then
				if wr='1' then --write
					tmp_ram(conv_integer(addr)) <= Din; 
				end if;
			end if;
	end process; 
	--Process #n...
	Dout<=(others=>'Z') when en='0' else tmp_ram(conv_integer(addr));--read 
end solve;